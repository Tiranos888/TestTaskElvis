
`timescale 1ns/1ps

// Main testbench module
module alu_tb;
logic clk;

// Test results counters
int passed_test_cnt;
int failed_test_cnt;

// Vector for test inputs 
logic [32:0] inputs_vector [100:0];

// Correct ALU output to check
logic [15:0] correct_alu_val = 16'h0000;

// Interface instantiation
alu_if alu_intf(clk);

// DUT instantiation using interface
alu16 dut (
//.clk(clk),
//.reset(alu_intf.reset),
.a(alu_intf.operand_a),
.b(alu_intf.operand_b),
.sel(alu_intf.opcode),
.mode(alu_intf.mode),
.Cin(alu_intf.carry_in),
.result(alu_intf.result),
.Cout(alu_intf.carry_out),
.nBo(), 
.nGo()
);

// Clock generation
initial begin
  clk = 0;
  forever #5 clk = ~clk;
end

// Test controller
initial begin
  initialize_test();
  run_tests();
  report_results();
  $finish;
end

// Helper tasks
task initialize_test();
  alu_intf.reset <= 1;
  alu_intf.operand_a <= 0;
  alu_intf.operand_b <= 0;
  alu_intf.opcode <= 0;
  alu_intf.carry_in <= 0;
  alu_intf.mode <= 0;
  #20;
  alu_intf.reset <= 0;
  $display("Test initialization completed");
endtask

task run_tests();
  test_add_operation();
  #20;
  test_sub_operation();
  #20;  
  test_inc_operation();
  #20;
  test_add_operation();
  #20;
  test_or_operation();
  #20;
endtask

// Individual test tasks
task test_add_operation();
  $display("Testing ADD operation...");
  alu_intf.opcode <= 4'b1001; // ADD
  alu_intf.mode <= 0;

  $readmemh("tests/add_operation_test", inputs_vector);
  
  for (int i = 0; i < 100; i++) begin
    if (inputs_vector[i] === 'x) break;

    {alu_intf.operand_a, alu_intf.operand_b, alu_intf.carry_in} = inputs_vector[i];

    @(posedge clk);
  end
  
endtask


task test_sub_operation();
  $display("Testing SUB operation...");
  alu_intf.opcode <= 4'b0110; // SUB
  alu_intf.mode <= 0;

  $readmemh("tests/sub_operation_test", inputs_vector);
  
  for (int i = 0; i < 100; i++) begin
    if (^inputs_vector[i] === 1'bX) break;

    {alu_intf.operand_a, alu_intf.operand_b, alu_intf.carry_in} <= inputs_vector[i];

    @(posedge clk);
  end

endtask


task test_inc_operation();
  $display("Testing INC operation...");
  alu_intf.opcode <= 4'b0011; // INC
  alu_intf.mode <= 0;

  $readmemh("tests/inc_operation_test", inputs_vector);
  
  for (int i = 0; i < 100; i++) begin
    if (^inputs_vector[i] === 1'bX) break;

    {alu_intf.operand_a, alu_intf.operand_b, alu_intf.carry_in} <= inputs_vector[i];

    @(posedge clk);
  end

endtask

task test_and_operation();
  $display("Testing AND operation...");
  alu_intf.opcode <= 4'b1100; // AND
  alu_intf.mode <= 1;

  $readmemh("tests/and_operation_test", inputs_vector);
  
  for (int i = 0; i < 100; i++) begin
    if (^inputs_vector[i] === 1'bX) break;

    {alu_intf.operand_a, alu_intf.operand_b, alu_intf.carry_in} <= inputs_vector[i];

    @(posedge clk);
  end
endtask


task test_or_operation();
  $display("Testing OR operation...");
  alu_intf.opcode <= 4'b1110; // OR
  alu_intf.mode <= 1;

  $readmemh("tests/or_operation_test", inputs_vector);
  
  for (int i = 0; i < 100; i++) begin
    if (^inputs_vector[i] === 1'bX) break;

    {alu_intf.operand_a, alu_intf.operand_b, alu_intf.carry_in} <= inputs_vector[i];

    @(posedge clk);
  end

endtask

// Results reporting
task report_results();
  $display("\n=== TEST SUMMARY ===");
  $display("All basic operations tested");
  $display("Testbench completed successfully");
  $display("%d tests passed", passed_test_cnt);
  $display("%d tests failed", failed_test_cnt);
endtask

function correct_alu_value(
    input [15:0] a,
    input [15:0] b,
    input [3:0]  opcode,
    input        carry_in
);

  case (opcode)
    4'b0000: correct_alu_value = a + b + carry_in;   // ADD
    4'b0001: correct_alu_value = a - b - carry_in;   // SUB
    4'b0101: correct_alu_value = {1'b0, a & b};      // AND
    4'b0110: correct_alu_value = {1'b0, a | b};      // OR
    4'b0111: correct_alu_value = {1'b0, a ^ b};      // XOR
    default: correct_alu_value = 17'hBAD1;
  endcase 
  
endfunction

always @(posedge clk) begin
  correct_alu_val = correct_alu_value(alu_intf.operand_a , alu_intf.operand_b , alu_intf.opcode , alu_intf.carry_in);

  if (alu_intf.result === correct_alu_val) begin
    $display("[PASS] A=%h B=%h res: %h", alu_intf.operand_a, alu_intf.operand_b, alu_intf.result);
    passed_test_cnt++;
  end else begin
    $display("[FAIL] A=%h B=%h exp=%h got=%h", alu_intf.operand_a, alu_intf.operand_b, correct_alu_val, alu_intf.result);
    failed_test_cnt++;
  end

end


// Additional monitoring
always @(posedge clk) begin
if (!alu_intf.reset) begin
  // Monitor can be extended here
  $display("Cycle: opcode=%h, a=%h, b=%h, result=%h, carry_out=%b",
            alu_intf.opcode, alu_intf.operand_a, 
            alu_intf.operand_b, alu_intf.result, alu_intf.carry_out);
end
end
endmodule